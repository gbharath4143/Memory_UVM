`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "memory.sv"

`include "common_mem.sv"
`include "txn_mem.sv"
`include "seq_mem.sv"
`include "interface_mem.sv"

`include "scoreboard_mem.sv"
`include "coverage_mem.sv"
`include "monitor_mem.sv"
`include "driver_mem.sv"
`include "sqr_mem.sv"
`include "agent_mem.sv"
`include "env_mem.sv"
`include "test_mem.sv"
`include "top_mem.sv"