class sqr_mem extends uvm_sequencer #(txn_mem);

  `uvm_component_utils(sqr_mem)

  `NEW_COMP

endclass